module multiplicator_nb()




endmodule 